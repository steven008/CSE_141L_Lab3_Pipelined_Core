library verilog;
use verilog.vl_types.all;
entity definitions_sv_unit is
end definitions_sv_unit;
