library verilog;
use verilog.vl_types.all;
entity miner_tb is
end miner_tb;
