library verilog;
use verilog.vl_types.all;
entity core_tb is
end core_tb;
