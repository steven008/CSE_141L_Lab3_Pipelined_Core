library verilog;
use verilog.vl_types.all;
entity cl_state_machine_sv_unit is
end cl_state_machine_sv_unit;
