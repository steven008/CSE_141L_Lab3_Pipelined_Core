library verilog;
use verilog.vl_types.all;
entity core_flattened_sv_unit is
end core_flattened_sv_unit;
