library verilog;
use verilog.vl_types.all;
entity core_sv_unit is
end core_sv_unit;
