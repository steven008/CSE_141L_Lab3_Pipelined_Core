library verilog;
use verilog.vl_types.all;
entity miner_tb_sv_unit is
end miner_tb_sv_unit;
