library verilog;
use verilog.vl_types.all;
entity cl_decode_sv_unit is
end cl_decode_sv_unit;
