library verilog;
use verilog.vl_types.all;
entity net_packet_logger_s_sv_unit is
end net_packet_logger_s_sv_unit;
