library verilog;
use verilog.vl_types.all;
entity instr_mem_sv_unit is
end instr_mem_sv_unit;
